
module TEST ( VDD, VSS, in, out );

    input VDD;
    input VSS;
    input in;
    output out;

endmodule
