
module TEST(
    input wire VDD,
    input wire VSS,
    input wire in,
    output wire out
);

endmodule
