
module TEST(
    inout wire B,
    inout wire D,
    inout wire G,
    inout wire S
);

endmodule
