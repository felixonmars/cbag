.PARAM

.SUBCKT nmos4_standard B D G S
.ENDS

.SUBCKT pmos4_standard B D G S
.ENDS

.SUBCKT cv_bus_term VDD VSS in<1> in<0> out
X3 VSS out in<1> VSS / nmos4_standard
X4 VDD out in<1> VDD / pmos4_standard l=90n nf=2 w=400n
XN VSS out in<0> VSS / nmos4_standard
XP VDD out in<0> VDD / pmos4_standard l=90n nf=2 w=400n
.ENDS

.SUBCKT TEST VDD VSS in<1> in<0> out
XINST VDD VSS in<1> in<0> out / cv_bus_term
.ENDS

