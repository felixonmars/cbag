
module TEST(
    input wire VDD,
    input wire VSS,
    input [1:0] wire in0,
    input [1:0] wire in1,
    output [1:0] wire out
);

endmodule
