.PARAM

.SUBCKT nmos4_standard B D G S
.ENDS

.SUBCKT pmos4_standard B D G S
.ENDS

.SUBCKT TEST VDD VSS in out
XN VSS out in VSS / nmos4_standard
XP VDD out in VDD / pmos4_standard l=90n nf=2 w=400n
.ENDS
