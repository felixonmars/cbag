.PARAM

.SUBCKT TEST B D G S
.ENDS

