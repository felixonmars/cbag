
module TEST(
    input wire VDD,
    input wire VSS,
    input [1:0] wire in,
    output wire out
);

endmodule
