
module TEST ( B, D, G, S );

    inout B;
    inout D;
    inout G;
    inout S;

endmodule
