
module TEST ( VDD, VSS, in, out );

    input VDD;
    input VSS;
    input [1:0] in;
    output out;

endmodule
