
module TEST ( VDD, VSS, in0, in1, out );

    input VDD;
    input VSS;
    input [1:0] in0;
    input [1:0] in1;
    output [1:0] out;

endmodule
