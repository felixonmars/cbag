.PARAM

.SUBCKT nmos4_standard B D G S
.ENDS

.SUBCKT pmos4_standard B D G S
.ENDS

.SUBCKT TEST VDD VSS in<1> in<0> out
XN<1> VSS out in<1> VSS / nmos4_standard
XN<0> VSS out in<0> VSS / nmos4_standard
XP<1> VDD out in<1> VDD / pmos4_standard l=90n nf=2 w=400n
XP<0> VDD out in<0> VDD / pmos4_standard l=90n nf=2 w=400n
.ENDS
